V1 1 0 5
R2 1 2 470
R3 0 2 330
.print dc v(2)
.dc
.end
